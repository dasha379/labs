module priority_encoder_4_tb;
  logic [3:0] data_i_tb;
  logic       data_val_i_tb;
  logic [3:0] data_left_o_tb;
  logic [3:0] data_right_o_tb;
  logic       data_val_o_tb;
  
  priority_encoder_4 DUT (
    .data_i      ( data_i_tb       ),
	 .data_val_i  ( data_val_i_tb   ),
	 .data_left_o ( data_left_o_tb  ),
	 .data_right_o( data_right_o_tb ),
	 .data_val_o  ( data_val_o_tb   )
  );
  
  task test
  (
    input [3:0] tdata,
	 input       tdata_val_i
  );
    logic [3:0] tdata_left, tdata_right;
	 logic tdata_val_o;
    
	 { data_i_tb, data_val_i_tb } = { tdata, tdata_val_i };
	 
	 #1ns;
	 
	 if (tdata_val_i == 0) 
		{ tdata_right, tdata_left, tdata_val_o } = { 4'b0, 4'b0, 1'b0 };
    else begin
      casez( tdata )
		  4'b1??? : tdata_left = 4'b1000;
		  4'b01?? : tdata_left = 4'b0100;
		  4'b001? : tdata_left = 4'b0010;
		  4'b0001 : tdata_left = 4'b0001;
		  default : tdata_left = 4'b0000;
	   endcase
			
		casez( tdata )
		  4'b1000 : tdata_right = 4'b1000;
		  4'b?100 : tdata_right = 4'b0100;
		  4'b??10 : tdata_right = 4'b0010;
	     4'b???1 : tdata_right = 4'b0001;
		  default : tdata_right = 4'b0000;
		endcase
		tdata_val_o = 1;
	 end
	 
	 if ( tdata_right != data_right_o_tb )  
	   $error("expected: %b, got: %b", tdata_right, data_right_o_tb);
    if ( tdata_left != data_left_o_tb )  
	   $error("expected: %b, got: %b", tdata_left, data_left_o_tb);
	 if ( tdata_val_o != data_val_o_tb )  
	   $error("expected: %b, got: %b", tdata_val_o, data_val_o_tb);
	 
  endtask
  
  initial begin
    test(4'b1111, 1);
	 test(4'b0000, 1);
	 test(4'b1111, 0);
	 test(4'b0000, 0);
	 
	 // test which covers all the cases without $random
	 for ( int i = 0; i < 15; i++ ) begin
		test(i, 1);
		test(i, 0);
	 end
    
	 // 5 random iterations
    for ( int i = 0; i < 5; i++ ) begin
	   data_i_tb = $urandom_range(15);
		data_val_i_tb = $urandom_range(1);
		test(data_i_tb, data_val_i_tb);
	 end
	 
	 $display("simulation is over, 0 errors");
	 $finish;
  end
  
endmodule